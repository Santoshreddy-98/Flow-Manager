jhwufhjwefn